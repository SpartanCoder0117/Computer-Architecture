Library ieee;
use ieee.std_logic_1164.all;
library lattice;
use lattice.componentes.all;

entity shiftRotate00 is 
port(
	clksl: in std_logic;
	enable: in std_logic;
	insl: in std_logic_vector(7 downto 0);
	sel: in std_logic_vector(3 downto 0);
	outsl: out std_logic_vector(7 downto 0)
	);
end shiftRotate00;

architecture shiftRotate0 of shiftRotate00 is 
signal sinsl: std_logic_vector(7 downto 0);
begin 
	psl: process(clksl)
	begin
		if (clksl'event and clksl = '1') then 
			case sel is
				when "0001" =>
					case enable is 
						when '0' => 
							outsl <= (others => '0');
							sinsl <= insl;
						when '1' => 
							sinsl(0) <= '0';--Desplazamiento derecha
							sinsl(7 downto 1) <= sinsl(6 downto 0);
							outsl <= sinsl;
					end case;
				when "0011" =>
					case enable is 
						when '0' => 
							outsl <= (others => '0');
							sinsl <= insl;
						when '1' => 
							sinsl(7) <= '0';--Desplazamiento izquierda
							sinsl(6 downto 0) <= sinsl(7 downto 1);
							outsl <= sinsl;
					end case;
				when "0111" =>
					case enable is 
						when '0' => 
							outsl <= (others => '0');
							sinsl <= insl;
						when '1' => 
							sinsl(0) <= sinsl(7);--Rotaci�n Izquierda
							sinsl(7 downto 1) <= sinsl(6 downto 0);
							outsl <= sinsl;
					end case;
				when "1111" =>
					case enable is 
						when '0' => 
							outsl <= (others => '0');
							sinsl <= insl;
						when '1' => 
							sinsl(7) <= sinsl(0);--Rotaci�n Izquierda
							sinsl(6 downto 0) <= sinsl(7 downto 1);
							outsl <= sinsl;
					end case;
				when others => null;
			end case;
		end if;
	end process psl;
end shiftRotate0; 