library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library lattice;
use lattice.components.all;

entity muxra00 is
	port();
end muxra00;

architecture muxra0 of muxra00 is
begin

end muxra0;
