library ieee;
library lattice;
use ieee.std_logic_1164.all;
use lattice.components.all;

entity pruebadis00 is
port(
	A,B,C,D : out std_logic
	);
end pruebadis00;

architecture pruebadis0 of pruebadis00 is
begin
	A <= '1';
B <= '1';C <= '1';
D <= '1';

end pruebadis0;